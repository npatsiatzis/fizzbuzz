library ieee;
	use ieee.std_logic_1164.all;
	use ieee.math_real.all;

package fizzbuzz_pkg is

end package fizzbuzz_pkg;